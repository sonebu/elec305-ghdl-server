saduadhadadaso